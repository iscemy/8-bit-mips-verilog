module adder (
    in1, in2, out
);
    
    
endmodule